package sv_mon_pkg;
    `include "../tb/models/sv_mon_logic/sram_mon.sv"
    `include "../tb/models/sv_mon_logic/utilization_mon.sv"
endpackage
