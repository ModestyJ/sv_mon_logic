package sv_mon_pkg;
    `include "sv_mon_logic/sram_mon.sv"
    `include "sv_mon_logic/utilization_mon.sv"
endpackage
