package sv_mon_pkg;
    `include "sram_mon.sv"
    `include "utilization_mon.sv"
endpackage
